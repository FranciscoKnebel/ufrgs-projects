--
-- Authors: Francisco Paiva Knebel
--				Gabriel Alexandre Zillmer
--
-- Universidade Federal do Rio Grande do Sul
-- Instituto de Inform�tica
-- Sistemas Digitais
-- Prof. Fernanda Lima Kastensmidt
--
-- Create Date:    17:04:14 05/14/2016 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity decimalTo7SEG is
	port (
		clk: 			in std_logic;
		bcd: 			in std_logic_vector(3 downto 0);
		segmented: 	out std_logic_vector(6 downto 0);
	);
end decimalTo7SEG;

architecture Behavioral of decimalTo7SEG is


begin
	if(clk'event AND clk = '1') then
		case bcd is
			segmented <= 	"0000001" when "0000", -- '0'
								"1001111" when "0001", -- '1'
								"0010010" when "0010", -- '2'
								"0000110" when "0011", -- '3'
								"1001100" when "0100", -- '4'
								"0100100" when "0101", -- '5'
								"0100000" when "0110", -- '6'
								"0001111" when "0111", -- '7'
								"0000000" when "1000", -- '8'
								"0000100" when "1001", -- '9'
								"0001000" when "1010", -- 'A'
								"1100000" when "1011", -- 'B'
								"0110001" when "1100", -- 'C'
								"1000010" when "1101", -- 'D'
								"0110000" when "1110", -- 'E'
								"0111000" when "1111", -- 'F'
								"1111111" when others;
		end case;
	end if;
end Behavioral;

